library verilog;
use verilog.vl_types.all;
entity fouroneMUX_vlg_vec_tst is
end fouroneMUX_vlg_vec_tst;
