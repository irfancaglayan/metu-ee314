library verilog;
use verilog.vl_types.all;
entity bcdCounter_vlg_vec_tst is
end bcdCounter_vlg_vec_tst;
